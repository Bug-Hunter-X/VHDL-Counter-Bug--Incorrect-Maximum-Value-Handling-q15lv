```vhdl
library ieee;
use ieee.std_logic_1164.all;

entity buggy_counter_fixed is
  port (
    clk : in std_logic;
    rst : in std_logic;
    count : out integer range 0 to 15
  );
end entity buggy_counter_fixed;

architecture behavioral of buggy_counter_fixed is
  signal internal_count : integer range 0 to 15 := 0;
begin
  process (clk, rst)
  begin
    if rst = '1' then
      internal_count <= 0;
    elsif rising_edge(clk) then
      case internal_count is
        when 15 => internal_count <= 0;
        when others => internal_count <= internal_count + 1;
      end case;
    end if;
  end process;
  count <= internal_count;
end architecture behavioral;
```